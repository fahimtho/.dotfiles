Vim�UnDo� �w�� Yh�z�ւ���3��v�5s_�Q�Vr��      	endmodule      	                      a�?s    _�                             ����                                                                                                                                                                                                                                                                                                                                                             a��     �                   5��                                                  �                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a�?`    �                   �               5��                                           �       5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                             a�?s     �               endmod5��                         �                      5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             a�?y    �               endmod:5��                         �                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��    �              �                 =module HELLO_WORLD(); // module doesn't have input or outputs     initial begin       $display("Hello World");   "    $finish; // stop the simulator     end   	endmodule5��                       	                   �       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             a��    �                endmodue5��                         �                      5��